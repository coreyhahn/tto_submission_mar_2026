`ifndef BYANG_PKG_VH
`define BYANG_PKG_VH

`define PRIME_BITS  256
`define OP_WIDTH    257
`define DELTA_WIDTH 10
`define NUM_ITERS   742
`define CTR_WIDTH   10
`define SECP256K1_P 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFC2F

`endif
